../../ADC_tb/systemVerilog/verilog.sv